module griffin_tb;

  // Parameters
  localparam N_BITS = 254;
  localparam PRIME_MODULUS = 254'h30644e72e131a029b85045b68181585d2833e84879b9709143e1f593f0000001;
  localparam BARRETT_R = 255'h54a47462623a04a7ab074a58680730147144852009e880ae620703a6be1de925;
  localparam STATE_SIZE = 3;
  localparam NUM_ROUNDS = 14;
  localparam CLK_PERIOD = 10; // 10ns clock period for 100 MHz clock
  
  // Inputs and Outputs
  reg clk;
  reg reset;
  reg enable;
  reg [N_BITS-1:0] inState [STATE_SIZE][13];
  wire [N_BITS-1:0] outState [STATE_SIZE][13];
  wire done;
    time start_time, end_time;
  // Test Vectors
  reg [N_BITS-1:0] testVector_1[STATE_SIZE*13];
  //reg [N_BITS-1:0] expectedVector [12][STATE_SIZE];
  
  // Instantiate the DUT
  griffin #(
    .N_BITS(N_BITS),
    .PRIME_MODULUS(PRIME_MODULUS),
    .BARRETT_R(BARRETT_R),
    .STATE_SIZE(STATE_SIZE),
    .NUM_ROUNDS(NUM_ROUNDS)
  ) dut (
    .clk(clk),
    .reset(reset),
    .enable(enable),
    .inState(inState),
    .outState(outState),
    .done(done)
  );
  
  // Clock generation
  initial begin
    clk = 0;
    forever #(CLK_PERIOD / 2) clk = ~clk;
  end

  // Test initialization and vector assignment
  initial begin
testVector_1[0] = 254'd19183296366840297261607075654228646741064326077950506146152119958439979864097;
testVector_1[1] = 254'd4145541186935938026593050205566893848843983243153598113321915732773859788351;
testVector_1[2] = 254'd10826373444134521561985703079771848275272288331843813040865871873516991765704;
testVector_1[3] = 254'd13059010918208593108840516037810737021500968883900878897087531485752054441776;
testVector_1[4] = 254'd18962205316629716089629550045781349996410263508838025262691497606025043166385;
testVector_1[5] = 254'd21690595958896654773242916386694403137299006628807566917516254018927139426768;
testVector_1[6] = 254'd5783661087944809595360845793696567520915671280836123294983292365757143229226;
testVector_1[7] = 254'd1469123457913188069101400702126786136560629096678798972410169925466448448424;
testVector_1[8] = 254'd12521300479215468644919198612302506167495523179877046350617389170802716379552;
testVector_1[9] = 254'd19473116388580141389032591771207874584755915878881382939147643628206069168648;
testVector_1[10] = 254'd11175019997888401711022850064888905062154712112269322475742785655155102117532;
testVector_1[11] = 254'd8652258866394102626161833837856845832809035066075201407074359983062031231888;
testVector_1[12] = 254'd5723934342698579566388545792479377786322174066748665471581872922956987607564;
testVector_1[13] = 254'd14441762024819145101563312900197271935433757243634442358857277566865458524453;
testVector_1[14] = 254'd5431803245163673298976842365073723058211043027681474475943116161740421237248;
testVector_1[15] = 254'd19520370316683093731719802927983557890256086175586465383333423001067383487871;
testVector_1[16] = 254'd13339616213015109345825002458705833605132322667027309331536391930989519148930;
testVector_1[17] = 254'd20436922409034520793965692692214297806629627496041500534582526246916461782729;
testVector_1[18] = 254'd18764907770179324051153353341835142085078612376154171345987645895951097747685;
testVector_1[19] = 254'd6873098683434528928059976161039078516855136952707773929571866369873510976375;
testVector_1[20] = 254'd10308958932719677747283778537406565112470406926683357228987760894100332292130;
testVector_1[21] = 254'd1249169345949784524964855429711449940529535943731343235391962195486771670400;
testVector_1[22] = 254'd3186635281795353972101562547598207898460383479097088651952210749978632276061;
testVector_1[23] = 254'd12218301402195486376443806165731614872580552908260829499993774131958041517833;
testVector_1[24] = 254'd2300294929772158011405127391373343360703354444240793700720222120249982333713;
testVector_1[25] = 254'd5809625220694393238157569615612389671746093850556705662627995764004041759810;
testVector_1[26] = 254'd18779125659766095679587997652319628327081884848497819919219193669738859198148;
testVector_1[27] = 254'd5957923925081643019715130710860620413793722037983904528875544661238317272402;
testVector_1[28] = 254'd1417765317980092617695561343387852538338397354720835260057582354060035953397;
testVector_1[29] = 254'd20341478657732359485015097777465126710742012188813049535518454386625878495223;
testVector_1[30] = 254'd14300997949432201924743277685599246443944405833844689704363257305644364039746;
testVector_1[31] = 254'd7071858593425000602801186179750089534735017278159141702530112743926480820156;
testVector_1[32] = 254'd590665616571927512988326133754589685197369799085150979574811949155772373156;
testVector_1[33] = 254'd11346740220691630857148898955135667519757521554470402151610280345499670357791;
testVector_1[34] = 254'd20061625505267518973076494615914930073089394071518635780390141135042462385112;
testVector_1[35] = 254'd13853530549069791879699142905485692307325268623244667738444995055667273881820;
testVector_1[36] = 254'd9316418872520697207326607613630008938336898439318906321463318135026215730167;
testVector_1[37] = 254'd1228118886911194995007031869401821156972588644036210345341629112411777043661;
testVector_1[38] = 254'd5755431680451793552524807876072280996525815020491463183965467442175681133236;

    // Reset and Initialize test
    reset = 1;
    enable = 0;
    #20 reset = 0;
    #10 enable = 1;

    // Capture the start time
    start_time = $time;

    // Begin test process
    for (int i = 0; i < 13; i++) begin
      for (int j = 0; j < STATE_SIZE; j++) begin
        inState[j][i] = testVector_1[3 * i + j];
      end
    end

    // Wait until computation completes
    wait (done);

    // Capture the end time
    end_time = $time;

    // Print elapsed time
    $display("Computation completed in %0t time units.", end_time - start_time);

    #100 $stop;
  end
  
endmodule



/*
Reference Input and Output:
Input: [FpBN254(0x2f9538bcb77a6521a0b7f22d254d119ac306ef4c22fb75c6850496297b8cf251), FpBN254(0x1b9440a8465faa450cb336897b6aa7c1286a6d9f8c3fa192f3f76b64456e3037), FpBN254(0x17ff4438ac3cb8f6d0a009045a33e993a02ee8518f6f1e0a047b25da4009c7ff)]
 Input: [FpBN254(0x0643f8f3395dc8b0e8b408b82b721443c297a678a824ae3f542250ad2067a1e2), FpBN254(0x1e708fe900637e529b30f06c1abe5fc67768d41f9f972e9d8bffeb5f13a1137a), FpBN254(0x2b0eb39bd5a78d5b7743f604a2d7471ca6d719534a49f43b7e554f75b259919f)]
 Input: [FpBN254(0x238bd30b6415b0fae9ec499dd256e395ede9ee198e93e316bfb808298d8bd8b8), FpBN254(0x0a269aa699f0231409d0b0dcf2f8cd23872f18fa3a97d8dc28a909925bb7bb33), FpBN254(0x152f0d09752dd2aac27ef40c7d374181dee3609591f10e21cac8d3b05685382f)]
 Input: [FpBN254(0x15f692f8bf4b01c16480c2bb92fabd0192029d3470fb2a6a4d4931da2d452f29), FpBN254(0x08a6ed4f0dc4d9165ee0cd491f601d775a3568f5ab8ad559b0f26543ce074773), FpBN254(0x0cec772704f61b6afc77770f4654bead5021e506484199f3856ca9373b2c9ff3)]
 Input: [FpBN254(0x0a8e568e0131308f7e47a7353730ad276c98e4ac8b7b27fb49011a2d5430efc2), FpBN254(0x0e9c4e07382362b8a86547257dddcee0301df49e3de9240686965d3bed70412b), FpBN254(0x05796e53a6db4f76a5b9eb9b0f448eaa548eef5d528663adc6aa35fc44dfbca9)]
 Input: [FpBN254(0x0cd736b196dee18fed80b42613b87e5aa8fde61dd3eaaa357e27bee426554980), FpBN254(0x2ae98af4f2fa443fd9903a861335626e32b43a6d395d5467b129fada065e7f37), FpBN254(0x1015ed96078108fb4e5d2c66e9b0b32c51e4d59d91e99793752161bf702a6ad4)]
 Input: [FpBN254(0x0f1bbcd632d94f034887987bad5e4677f2119a5f3ef66ef3cddfef025db76ab9), FpBN254(0x26b52eeb58bc2eec8faf95345dc3fe28ce635a35b69805ef0706068f791cfe64), FpBN254(0x0dad286152db9007f2912bfaadbd633a6e65235419de5f91ff7f8f749f6b7885)]
 Input: [FpBN254(0x0dd552e6b63d0d6bea182a18cd34dc8813e5c702c43f43f448cb8e9636e32398), FpBN254(0x05ab412ab0e71702afc1f059d0e64788d0665874d9e5a1b23f0f76a059433172), FpBN254(0x13ae40e7a84ec05f8a59b016996274f516be60ae3c843f8ce1128ac275d11f68)]
 Input: [FpBN254(0x299810a4f8e9ea074f046eb7e341616db10cd5772a8ad6c63fe8c0b8fabfdc1a), FpBN254(0x077a46db19166d5bc8290b3ff0873e9776cc7c79190d5ae9a0bb2b8c9c1180f5), FpBN254(0x0b6fa2da4c29d70e7ca729fac9eeba578f0fbb5defb5589a83c8caa0f21de5b0)]
 Input: [FpBN254(0x097efb3ae35c794b4cef6c9b655260f499bc04fe0d76ca1ede93c3d9bf6920d3), FpBN254(0x172c42f2ae1873010033b0af011b45774393b21c7331859ad80a60f0ac930aba), FpBN254(0x03ead04ff6edb25fe8d5736f961453720a3ea1b73651cc83e109de2054d71320)]
 Input: [FpBN254(0x068938c1eb701d63482631ff5dab1f97cb621d2450f4ade828adefeeca99c0d9), FpBN254(0x28d9a072260d40a5444b75cca31ace80ddc6fb11abbc8b296c87435d420f1429), FpBN254(0x26f04d3da39892de8ac039450b399b160364f4ba2d1da96f34749b582fa301fb)]
 Input: [FpBN254(0x1dc5f3db74d372b7053efb312b99ebc078d6088c71e06b4014c62953339e8c9b), FpBN254(0x18553423819d5baf5f3478534eb2e7fb8502c240c86e505454799b687fb72ef6), FpBN254(0x0d6fa16776eaf7958af9da184929234a994651fe93c140da977eab55f260d5c9)]
 Input: [FpBN254(0x1b18ace654e632fce7a9876dcab29239ce4963f816ff0610b619dd7642c64624), FpBN254(0x148bde7b710dca18f23e49dc1f1d44504945455ede41c9c5dd1f56409632c0c0), FpBN254(0x1d81db2750a71d442bf370afd26b7cfd4a902c5d9c0876ec8e03387c225a6887)]
 Permuted Output: [FpBN254(0x2fbfccf712dc3a8a062742550c7f4771e52fdc2f328da38fec4191d7db78969d), FpBN254(0x10f2a33cda7417b91e7e218dc68ee3ef4b6238520d18708ca1bdcbd1636385db), FpBN254(0x2e1ab9e38ba3f321df26fa05eec12ca6cc04b927759d22bbe7c958c2c4a358b0)]
 Permuted Output: [FpBN254(0x1da8c4b90095c05e715cc5459a487842b96d391fd7de81901ec5167b665f2a22), FpBN254(0x2ec594e97ae6e8f467208e84cad2177f3900faa7b4fc0089f5cd23375a733624), FpBN254(0x1767f05ca3b66c587b0b5fb7e634f5015a72b0fb27ddacbd9b76ccb97476bf9f)]
 Permuted Output: [FpBN254(0x01b025068a65dd4cbd816e70edead55ae484fbf6f4ef61e59d13ad65f797addb), FpBN254(0x28c703198cba778413db40e232e28d0ab16bd4d034fba88597bdb5dadd66f184), FpBN254(0x0b0eeac5e4759bf9eb1c754de734fcb87f08fa24fb39edd988875d8b10a9e4f1)]
 Permuted Output: [FpBN254(0x1c29de1a356ba9956af95fce11e91bf03826ebf8943d82636265ad71409c1d3b), FpBN254(0x278d05c91b7fc7fe16608eb444a4e5220449f9303d92060f1ed74779f6fde2dc), FpBN254(0x293ef812d787525c20556b44c8ea49dcb3474c6d38e2332b5049999c7661eacd)]
 Permuted Output: [FpBN254(0x096648192d426a46f4a30695ab07c4146dbae1014f2232dced92a80a0d8ba6a0), FpBN254(0x2dc6fea2bdb3156f748b17c15b13a8a091dd9171dfb4d8be472daa515a4bd2e2), FpBN254(0x22ba6b007d2ad0bb7c3649eadf8b9e41020ac0da6d4d75240d405ecba8eeb1ff)]
 Permuted Output: [FpBN254(0x2c40f4dc18a0d38a45d5801160063f89f60ac2af11475237176c966e042720a3), FpBN254(0x045cd2d97d277dfc7a71489bf9a35e13748f7522cf864d28607ed057504b2602), FpBN254(0x1a0853e09ddb99f52c2895965b25ae16ba41b542601297d35dd67fd429ed4022)]
 Permuted Output: [FpBN254(0x300def7a3e6f080cdb0a2f0e333d76966dfefc1c42e4162b75f9ce4f9199d4ac), FpBN254(0x2d06ce54f576970e187ae8424b5d080301f5370339017f1d2d99c5720b0a4e92), FpBN254(0x05cde8a7a5c51a80d9ee6cf30a48359fe0c28aa182cd1d47c290729c0541f34e)]
 Permuted Output: [FpBN254(0x16eedc2349f8c44bc54f6ad0f92cef8947926372c067461abca740fedc8b52af), FpBN254(0x19ff4c037c9d11ce4a9a14950c851a9c5f44c3b20ed08025377bf019b9df281b), FpBN254(0x28eea1d9bbe75f5a6f0b432c545095906c87955748eca5f5bc4de8c54969b3f8)]
 Permuted Output: [FpBN254(0x0bf747c6db17b67b393a8a8a4a0e3e47dfcdba588001168403e9ba3f827e06fc), FpBN254(0x1f428fac6587d07ee7298d06390e53539b2e6926660605ab4e9544a6d6c4d1f3), FpBN254(0x240b5c1e21e070a3fcdd7cd2a964551d47e54a56847172e639b09e48ff6ceed5)]
 Permuted Output: [FpBN254(0x1f15e76452be89c384650d8e6d0c75b135fe406a1119e99e2086e550bc66b4cd), FpBN254(0x066fe346c642fcc7ab0a66229cce1492e01076753706c2acbb0d9b181494d202), FpBN254(0x26c3d794536367db0d534b0ef74802ba231b693a153c0fede8c9a59690374a9e)]
 Permuted Output: [FpBN254(0x04c971e4fbbf96ca3f12e9af21be4c2d88ee94fe9c15e9ff7a51b7ae4ced5723), FpBN254(0x1570114956e966250b6352009b376ebf524ccc6f865543533148486044c9afef), FpBN254(0x158a5b4f2c41e9fb9ae86307c6c58a20ee19850751d5d1ded0b1148238af9984)]
 Permuted Output: [FpBN254(0x21ec76292069dc6b196a97814fc77e4fa09869399cff347bd0396281ea1d3141), FpBN254(0x1e4620d096c8c28e45afefd87609dc6c5339e9ae3342f60a32030c642ba8c5e0), FpBN254(0x212fb94e1a265aa9b75bb9e4101f12ba11b49ab51af2935602bc2bdfd6d61915)]
 Permuted Output: [FpBN254(0x23a9bba6c60e6ac1489892c51048a67884fbf6ee7cae889d91db83e748935481), FpBN254(0x09991d896814dd54c3211634fe9b03b2e12f3907bb1f5b2856f1fa5ea218fa2e), FpBN254(0x16afbfc998efba58af670eb9aa636d08e18eb74cbe52a5a46379dda68ee835d3)]

*/