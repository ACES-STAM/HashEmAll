/*
Reference input and output(in decimal):
Permutation - Input: [7, 5, 0]
Permutation - Output: [12360106593270449844061412657301362366573579256583003766552363058581964117186, 571281065699991603834232145226702411332243584689159097661681181035646779147, 5827211446942541137487801220137246525465448099690109106563675347241842025991]
Permutation - Input: [10917901770635866436075026016659080286184149548927087489003364430639471220657, 15093033869696199585334196511061284287566496673224764407232042360381732406822, 0]
Permutation - Output: [9015251630996607203618061446630382221872903244076542510604305929244679444419, 15879859090627996012910608502246148008395297925036347252664944182065690596621, 18560181493604561726790764277907035345951571022315713369595937606897153822615]
Permutation - Input: [21739712095178135048191546448963631920285197592697942392244793527788985886301, 8858283708315735321250403702432677061468885569337168495636056784571574406448, 0]
Permutation - Output: [18329931618415610668643634474014011335241935075190086161442182803215507500299, 2149369278479666633097953201825936302312307642502164003213072662610116947450, 1803625172765819007712227852553682169356933782067426899770176074186941360527]
Permutation - Input: [15647695940089500251678240681748798303434417819422794141800595102470224949797, 18478792838189852650095108189496860401827254585568628862804027353559861163985, 0]
Permutation - Output: [20486877510231618053066305798476308324104477256085821770670638367672575655972, 8506186614711587338271697025571522047350453599120149045311718895163873227158, 19331295163941894760549037142871984830693281730919883221311891988423964809664]
Permutation - Input: [19900524514612089806276604711837690453215070955832409975167381678422194897905, 1236606864354083188154591020243375615684840709595277385538149191988208506003, 0]
Permutation - Output: [15009369781091431499304070154912425359963382052464747391162946304596761648983, 17956993152787252927978581752944873836913007540812860576695818296736105965895, 20851007939158033029485606678152121739648672092401282804037817306968291308858]        
Permutation - Input: [20767081487668653306571970702982492773897412604424936666057505328864346471759, 5272159900800745762041740216767697914529812765717334033541487238715296148735, 0]
Permutation - Output: [20391782752823351916950710951584738593182576402115041728038492224577649332407, 21883934090929647172947679351779169281356816682663455117570507161160307800396, 17973598412196279653593606919328301226782415401620279915007894720105912403962]        
Permutation - Input: [9375207379161327853834308035010312852168568912774835926127390746572711653001, 18215294625592889596659303014994370765104507296543683038994134854673879109294, 0]
Permutation - Output: [19889201785444021530172424054140421604460547437976494848908655224396167553691, 5044671079490109332583090548905605047119878548832898313009479887641901576083, 1929933356026833760244198349596534755426312920563985950859654429696970425113]
Permutation - Input: [10442286909081447267778762487686955053420267485148173562551203049360125464309, 16414624291395617007545606219325363297485841380931547081432204698622829918059, 0]
Permutation - Output: [586931882465379973006570884560276388695335080962126786585334541594909638309, 10605590130054669982856577385566522123140177003613674829813146832297847874258, 12307656769483557841410822449766043069022688507182348556505429197287396560879]
Permutation - Input: [18837118988058782052907318170698452279560628312810076072342995247067701518258, 16705760111171223003951385386167643144584727294835379247504400984470192160688, 0]
Permutation - Output: [16596004394661610479122068598376906184305117752428815886081358879375591503791, 6741503635933551527107418409987439049104817672199007442045349756558814744489, 5558053279613392977281211721557313500134533314227567752367454852364877174955]
Permutation - Input: [5668094874103265696334551985640714133195387871229321113793698399566639512531, 5741960809815986019555904263416509216658722978137227432436430694971609592605, 0]
Permutation - Output: [20312383426545192611004893133874574752818372414797828357655346399368693793943, 4708829991803901504383743674115403649678177031808853369532565347040106996692, 12909228403971079314776936413852458583437435034074953780080402131569686453688]
Permutation - Input: [6087197294869114683777430443143440645720269033823964295565433563153171048140, 613784097092740180855052074166703620398728665939444412094895167860409273165, 0]
Permutation - Output: [11353501954590241139520956562143277668647705157009295084684059358521690511653, 4703085232975642147986339022696158401290520001257460041363588534276401671182, 8043069950384460949795636221448758395401471276227686134376467133418819805160]
Permutation - Input: [15456325924657491730148759865200832894571452057020814710844324085824832797932, 12266559940464367019075897177603685313945104910251119269749009731576014557555, 0]
Permutation - Output: [16682507527068287853940624795376103653397356963636959815185582131350975175551, 18897809649774000760636094983135481539778060017780735747681166112838742221360, 5754732557433427612157190016632686976712472482376761166933319574849245848156]
Permutation - Input: [1485130523526814394494219916554092458724911195344785758817920831066365205568, 10649320480001284802605218039042849994260571124891269262416666201188633701405, 0]
Permutation - Output: [19353883476287036883511347389610418528563609215800791665646647733738502746470, 12087580417395704682787375847542600002016002977387736481424707135723089961574, 1756968207129097057878199120117796069656823716921756986264483855510770593187]
*/


module tb_rcPermutation;

// Parameters
localparam STATE_SIZE = 3;
localparam N_BITS = 254;
localparam PRIME_MODULUS = 254'h30644e72e131a029b85045b68181585d2833e84879b9709143e1f593f0000001;
localparam BARRETT_R = 255'h54a47462623a04a7ab074a58680730147144852009e880ae620703a6be1de925;

// Testbench signals
logic clk, reset, enable;
  logic [N_BITS-1:0] inState[STATE_SIZE][13];
  logic [N_BITS-1:0] outState[STATE_SIZE][13];
logic done;
  logic [N_BITS-1:0] testVector1[STATE_SIZE*13];
// Time measurement variables
time start_time, end_time;

// DUT instance
rcPermutation #(
    .STATE_SIZE(STATE_SIZE),
    .N_BITS(N_BITS),
    .PRIME_MODULUS(PRIME_MODULUS),
    .BARRETT_R(BARRETT_R)
) dut (
    .clk(clk),
    .reset(reset),
    .enable(enable),
    .inState(inState),
    .outState(outState),
    .done(done)
);

// Clock generation
initial clk = 0;
always #5 clk = ~clk; // 10ns period

// Testbench variables
integer i;

initial begin
testVector1[0] = 254'd7;
testVector1[1] = 254'd5;
testVector1[2] = 254'd0;
testVector1[3] = 254'd10917901770635866436075026016659080286184149548927087489003364430639471220657;
testVector1[4] = 254'd15093033869696199585334196511061284287566496673224764407232042360381732406822;
testVector1[5] = 254'd0;
testVector1[6] = 254'd21739712095178135048191546448963631920285197592697942392244793527788985886301;
testVector1[7] = 254'd8858283708315735321250403702432677061468885569337168495636056784571574406448;
testVector1[8] = 254'd0;
testVector1[9] = 254'd15647695940089500251678240681748798303434417819422794141800595102470224949797;
testVector1[10] = 254'd18478792838189852650095108189496860401827254585568628862804027353559861163985;
testVector1[11] = 254'd0;
testVector1[12] = 254'd19900524514612089806276604711837690453215070955832409975167381678422194897905;
testVector1[13] = 254'd1236606864354083188154591020243375615684840709595277385538149191988208506003;
testVector1[14] = 254'd0;
testVector1[15] = 254'd20767081487668653306571970702982492773897412604424936666057505328864346471759;
testVector1[16] = 254'd5272159900800745762041740216767697914529812765717334033541487238715296148735;
testVector1[17] = 254'd0;
testVector1[18] = 254'd9375207379161327853834308035010312852168568912774835926127390746572711653001;
testVector1[19] = 254'd18215294625592889596659303014994370765104507296543683038994134854673879109294;
testVector1[20] = 254'd0;
testVector1[21] = 254'd10442286909081447267778762487686955053420267485148173562551203049360125464309;
testVector1[22] = 254'd16414624291395617007545606219325363297485841380931547081432204698622829918059;
testVector1[23] = 254'd0;
testVector1[24] = 254'd18837118988058782052907318170698452279560628312810076072342995247067701518258;
testVector1[25] = 254'd16705760111171223003951385386167643144584727294835379247504400984470192160688;
testVector1[26] = 254'd0;
testVector1[27] = 254'd5668094874103265696334551985640714133195387871229321113793698399566639512531;
testVector1[28] = 254'd5741960809815986019555904263416509216658722978137227432436430694971609592605;
testVector1[29] = 254'd0;
testVector1[30] = 254'd6087197294869114683777430443143440645720269033823964295565433563153171048140;
testVector1[31] = 254'd613784097092740180855052074166703620398728665939444412094895167860409273165;
testVector1[32] = 254'd0;
testVector1[33] = 254'd15456325924657491730148759865200832894571452057020814710844324085824832797932;
testVector1[34] = 254'd12266559940464367019075897177603685313945104910251119269749009731576014557555;
testVector1[35] = 254'd0;
testVector1[36] = 254'd1485130523526814394494219916554092458724911195344785758817920831066365205568;
testVector1[37] = 254'd10649320480001284802605218039042849994260571124891269262416666201188633701405;
testVector1[38] = 254'd0;
    $dumpfile("tb_rc_permutation.vcd");
  $dumpvars(0, tb_rcPermutation);

    // Initialize inputs
    reset = 1;
    enable = 0;

    // Apply reset
    #20;
    reset = 0;

    // Apply input stimulus
    #10;
    enable = 1;
    start_time = $time; // Record the start time
	
  for(int i = 0; i < 13;i++) begin
    for(int j = 0; j < STATE_SIZE; j++) begin
      inState[j][i] = testVector1[3*i+j];
    end
  end

    // Wait for the computation to complete
    wait (done);
    end_time = $time; // Record the end time
    $display("Computation completed.");
    $display("Time elapsed: %0t ns", end_time - start_time);

//     // Display the outputs
//     for (i = 0; i < STATE_SIZE; i++) begin
//         $display("outState[%0d] = %d", i, outState[i]);
//     end

    // Finish simulation
    #20;
    $stop;
end

endmodule
