`include "affine_3.sv"
`include "galois_add_three.sv"
`include "griffinPi.sv"
`include "galois_mult_barrett_sync.sv"
`include "mult_256_sync.sv"
`include "galois_pow_5.sv"
`include "galois_pow_dinv.sv"
`include "galois_mult_254.sv"
`include "Li.sv"
`include "nonlinear.sv"
`include "griffinPi.sv"
`include "griffin.sv"
`include "griffin_top.sv"