module tb_rescuePrime;

    // Parameters
    parameter N_BITS = 254;
    parameter PRIME_MODULUS = 254'h30644e72e131a029b85045b68181585d2833e84879b9709143e1f593f0000001;
    parameter BARRETT_R = 255'h54a47462623a04a7ab074a58680730147144852009e880ae620703a6be1de925;
    parameter STATE_SIZE = 3;
    parameter NUM_ROUNDS = 14;

    // Inputs
  reg [N_BITS-1:0] inState[STATE_SIZE][13];
    reg clk, enable, reset;

    // Outputs
  wire [N_BITS-1:0] outState[STATE_SIZE][13];
    wire done;
  logic [N_BITS-1:0] testVector[STATE_SIZE][13];
    // Instantiate the Unit Under Test (UUT)
    rescuePrime #(
        .N_BITS(N_BITS),
        .PRIME_MODULUS(PRIME_MODULUS),
        .BARRETT_R(BARRETT_R),
        .STATE_SIZE(STATE_SIZE),
        .NUM_ROUNDS(NUM_ROUNDS)
    ) uut (
        .inState(inState),
        .clk(clk),
        .enable(enable),
        .reset(reset),
        .outState(outState),
        .done(done)
    );

    // Clock generation
    initial clk = 0;
    always #5 clk = ~clk; // 10ns clock period

    // Stimulus
    initial begin
      $dumpfile("tb_rescuePrime.vcd");
      $dumpvars(0,tb_rescuePrime);
      testVector[0][0] = 254'd14382792074241024997102314384864298448063038247118480295047980188218088024987;
testVector[1][0] = 254'd21619987514702361662314720973711248711016328709023131247678554389934151420184;
testVector[2][0] = 254'd10065590997828011040291204352866097011201627908723464555802919279363754034169;
testVector[0][1] = 254'd17734352908045968852542945006759484205357847114740036386697763092459420498316;
testVector[1][1] = 254'd4690971412162320167945543024621611097976420827463383157122600400956925749207;
testVector[2][1] = 254'd9886272910761008459304253768797029799095306207839584202105231568503736799021;
testVector[0][2] = 254'd13486087979922436734101767003175437605600004034144364183353517140425161957322;
testVector[1][2] = 254'd15321816511580413002581308548543062000502493055519160857823621566964293091525;
testVector[2][2] = 254'd10597819961622776181390933356886031186819118312074379738693313433048259837361;
testVector[0][3] = 254'd3347263821600633527587740815985119000867919685776812063941189462221044055183;
testVector[1][3] = 254'd17976989309370486445429994952948247398255173709069914357676367845941743157530;
testVector[2][3] = 254'd11882134319984635335448141337028653003061352540707560597420442269748410309559;
testVector[0][4] = 254'd4361161864957802791584289739027758593146224150365766230348751378074567607842;
testVector[1][4] = 254'd12588831239024800279263721074186439615072102032728726216358535481403719726315;
testVector[2][4] = 254'd4163171600349492766266770004030570932551331826008978556995471574999973748546;
testVector[0][5] = 254'd13386196442948941201469676743141613691966941599214589598811123044573874815201;
testVector[1][5] = 254'd1147794990119410545625486976098858521234372068158482743841405529016952085271;
testVector[2][5] = 254'd20544258417884931681784146763280741557245648946236085635016737681961252787423;
testVector[0][6] = 254'd21403346990480878164287574976876784314947697587793871276212864925525834310013;
testVector[1][6] = 254'd14494371062046996377289962672658981121418045128890264075698691636074632476887;
testVector[2][6] = 254'd8816725860368372832583417987326658859751460602834936943070409823227210346067;
testVector[0][7] = 254'd5408584758667275474657459131420364374174747814896427340569886620587441219984;
testVector[1][7] = 254'd2398333394068243698189867245095528906489966064337321202928374639523035491082;
testVector[2][7] = 254'd17500708409707160164627368599825255002443724037115348993857836957605782475090;
testVector[0][8] = 254'd16820749526648346293356580992879592944502695957256438906149546411033219909252;
testVector[1][8] = 254'd17122086957655602137863741210329109315746423829003408926514332645103392764524;
testVector[2][8] = 254'd6689723944572337753138998383030624001009025622982851528872124630412083642253;
testVector[0][9] = 254'd6739819659053004844804608174576234407684495701043719715738018042678209135019;
testVector[1][9] = 254'd6487053258539889236836245528154298753131398759041426552001721173361744991045;
testVector[2][9] = 254'd8025412158605764034549980014456195968561855255273219276564309538788122480589;
testVector[0][10] = 254'd16734270622016618569600350917511627223164215105684433058397386875712496084761;
testVector[1][10] = 254'd21703250629052661482132067997598192199186976879399629279179459640402326243156;
testVector[2][10] = 254'd15393393828098230375066776286708715147701574890752213952943948745029835920483;
testVector[0][11] = 254'd4898928435969928282861794631911461540334938483280829669979147235048858108061;
testVector[1][11] = 254'd6242436518257294969600187942885620955900763187715870624850722326482609678685;
testVector[2][11] = 254'd15745885816229262717866944811284678430276183172638127391170027595980990619074;
testVector[0][12] = 254'd8708236930035547068445640451045807354234938758332712489026683032949678462293;
testVector[1][12] = 254'd11059343321715678319110373097325574374321963111813502841103361680682958078937;
testVector[2][12] = 254'd18515684859878303533458471264829859861386063584672169285773260112511296923332;
        // Initialize inputs
        reset = 1;
        enable = 0;
        // Reset the module
        #10 reset = 0;
        enable = 1;
      for (int i = 0; i < 13; i++) begin
        inState[0][i] = testVector[0][i];
        inState[1][i] = testVector[1][i];
        inState[2][i] = testVector[2][i];
      end
      #10 enable = 0;
        // Wait for the module to complete
        wait (done);
//       for(int i = 0; i < 13; i++) begin
//         for (int j = 0; j < 13; j ++) begin
        	
//           $display("outState[%1d][%1d] = %h", j, i, outState[j][i]);
//         end
//       end
        // Display output
        // End simulation
        #200 $stop;
    end

endmodule
