/*
Reference Input and Output(in hex):
Input: [FpBN254(0x2f9538bcb77a6521a0b7f22d254d119ac306ef4c22fb75c6850496297b8cf251), FpBN254(0x1b9440a8465faa450cb336897b6aa7c1286a6d9f8c3fa192f3f76b64456e3037), FpBN254(0x17ff4438ac3cb8f6d0a009045a33e993a02ee8518f6f1e0a047b25da4009c7ff)]
 Input: [FpBN254(0x0643f8f3395dc8b0e8b408b82b721443c297a678a824ae3f542250ad2067a1e2), FpBN254(0x1e708fe900637e529b30f06c1abe5fc67768d41f9f972e9d8bffeb5f13a1137a), FpBN254(0x2b0eb39bd5a78d5b7743f604a2d7471ca6d719534a49f43b7e554f75b259919f)]
 Input: [FpBN254(0x238bd30b6415b0fae9ec499dd256e395ede9ee198e93e316bfb808298d8bd8b8), FpBN254(0x0a269aa699f0231409d0b0dcf2f8cd23872f18fa3a97d8dc28a909925bb7bb33), FpBN254(0x152f0d09752dd2aac27ef40c7d374181dee3609591f10e21cac8d3b05685382f)]
 Input: [FpBN254(0x15f692f8bf4b01c16480c2bb92fabd0192029d3470fb2a6a4d4931da2d452f29), FpBN254(0x08a6ed4f0dc4d9165ee0cd491f601d775a3568f5ab8ad559b0f26543ce074773), FpBN254(0x0cec772704f61b6afc77770f4654bead5021e506484199f3856ca9373b2c9ff3)]
 Input: [FpBN254(0x0a8e568e0131308f7e47a7353730ad276c98e4ac8b7b27fb49011a2d5430efc2), FpBN254(0x0e9c4e07382362b8a86547257dddcee0301df49e3de9240686965d3bed70412b), FpBN254(0x05796e53a6db4f76a5b9eb9b0f448eaa548eef5d528663adc6aa35fc44dfbca9)]
 Input: [FpBN254(0x0cd736b196dee18fed80b42613b87e5aa8fde61dd3eaaa357e27bee426554980), FpBN254(0x2ae98af4f2fa443fd9903a861335626e32b43a6d395d5467b129fada065e7f37), FpBN254(0x1015ed96078108fb4e5d2c66e9b0b32c51e4d59d91e99793752161bf702a6ad4)]
 Input: [FpBN254(0x0f1bbcd632d94f034887987bad5e4677f2119a5f3ef66ef3cddfef025db76ab9), FpBN254(0x26b52eeb58bc2eec8faf95345dc3fe28ce635a35b69805ef0706068f791cfe64), FpBN254(0x0dad286152db9007f2912bfaadbd633a6e65235419de5f91ff7f8f749f6b7885)]
 Input: [FpBN254(0x0dd552e6b63d0d6bea182a18cd34dc8813e5c702c43f43f448cb8e9636e32398), FpBN254(0x05ab412ab0e71702afc1f059d0e64788d0665874d9e5a1b23f0f76a059433172), FpBN254(0x13ae40e7a84ec05f8a59b016996274f516be60ae3c843f8ce1128ac275d11f68)]
 Input: [FpBN254(0x299810a4f8e9ea074f046eb7e341616db10cd5772a8ad6c63fe8c0b8fabfdc1a), FpBN254(0x077a46db19166d5bc8290b3ff0873e9776cc7c79190d5ae9a0bb2b8c9c1180f5), FpBN254(0x0b6fa2da4c29d70e7ca729fac9eeba578f0fbb5defb5589a83c8caa0f21de5b0)]
 Input: [FpBN254(0x097efb3ae35c794b4cef6c9b655260f499bc04fe0d76ca1ede93c3d9bf6920d3), FpBN254(0x172c42f2ae1873010033b0af011b45774393b21c7331859ad80a60f0ac930aba), FpBN254(0x03ead04ff6edb25fe8d5736f961453720a3ea1b73651cc83e109de2054d71320)]
 Input: [FpBN254(0x068938c1eb701d63482631ff5dab1f97cb621d2450f4ade828adefeeca99c0d9), FpBN254(0x28d9a072260d40a5444b75cca31ace80ddc6fb11abbc8b296c87435d420f1429), FpBN254(0x26f04d3da39892de8ac039450b399b160364f4ba2d1da96f34749b582fa301fb)]
 Input: [FpBN254(0x1dc5f3db74d372b7053efb312b99ebc078d6088c71e06b4014c62953339e8c9b), FpBN254(0x18553423819d5baf5f3478534eb2e7fb8502c240c86e505454799b687fb72ef6), FpBN254(0x0d6fa16776eaf7958af9da184929234a994651fe93c140da977eab55f260d5c9)]
 Input: [FpBN254(0x1b18ace654e632fce7a9876dcab29239ce4963f816ff0610b619dd7642c64624), FpBN254(0x148bde7b710dca18f23e49dc1f1d44504945455ede41c9c5dd1f56409632c0c0), FpBN254(0x1d81db2750a71d442bf370afd26b7cfd4a902c5d9c0876ec8e03387c225a6887)]
 Permuted Output: [FpBN254(0x2fbfccf712dc3a8a062742550c7f4771e52fdc2f328da38fec4191d7db78969d), FpBN254(0x10f2a33cda7417b91e7e218dc68ee3ef4b6238520d18708ca1bdcbd1636385db), FpBN254(0x2e1ab9e38ba3f321df26fa05eec12ca6cc04b927759d22bbe7c958c2c4a358b0)]
 Permuted Output: [FpBN254(0x1da8c4b90095c05e715cc5459a487842b96d391fd7de81901ec5167b665f2a22), FpBN254(0x2ec594e97ae6e8f467208e84cad2177f3900faa7b4fc0089f5cd23375a733624), FpBN254(0x1767f05ca3b66c587b0b5fb7e634f5015a72b0fb27ddacbd9b76ccb97476bf9f)]
 Permuted Output: [FpBN254(0x01b025068a65dd4cbd816e70edead55ae484fbf6f4ef61e59d13ad65f797addb), FpBN254(0x28c703198cba778413db40e232e28d0ab16bd4d034fba88597bdb5dadd66f184), FpBN254(0x0b0eeac5e4759bf9eb1c754de734fcb87f08fa24fb39edd988875d8b10a9e4f1)]
 Permuted Output: [FpBN254(0x1c29de1a356ba9956af95fce11e91bf03826ebf8943d82636265ad71409c1d3b), FpBN254(0x278d05c91b7fc7fe16608eb444a4e5220449f9303d92060f1ed74779f6fde2dc), FpBN254(0x293ef812d787525c20556b44c8ea49dcb3474c6d38e2332b5049999c7661eacd)]
 Permuted Output: [FpBN254(0x096648192d426a46f4a30695ab07c4146dbae1014f2232dced92a80a0d8ba6a0), FpBN254(0x2dc6fea2bdb3156f748b17c15b13a8a091dd9171dfb4d8be472daa515a4bd2e2), FpBN254(0x22ba6b007d2ad0bb7c3649eadf8b9e41020ac0da6d4d75240d405ecba8eeb1ff)]
 Permuted Output: [FpBN254(0x2c40f4dc18a0d38a45d5801160063f89f60ac2af11475237176c966e042720a3), FpBN254(0x045cd2d97d277dfc7a71489bf9a35e13748f7522cf864d28607ed057504b2602), FpBN254(0x1a0853e09ddb99f52c2895965b25ae16ba41b542601297d35dd67fd429ed4022)]
 Permuted Output: [FpBN254(0x300def7a3e6f080cdb0a2f0e333d76966dfefc1c42e4162b75f9ce4f9199d4ac), FpBN254(0x2d06ce54f576970e187ae8424b5d080301f5370339017f1d2d99c5720b0a4e92), FpBN254(0x05cde8a7a5c51a80d9ee6cf30a48359fe0c28aa182cd1d47c290729c0541f34e)]
 Permuted Output: [FpBN254(0x16eedc2349f8c44bc54f6ad0f92cef8947926372c067461abca740fedc8b52af), FpBN254(0x19ff4c037c9d11ce4a9a14950c851a9c5f44c3b20ed08025377bf019b9df281b), FpBN254(0x28eea1d9bbe75f5a6f0b432c545095906c87955748eca5f5bc4de8c54969b3f8)]
 Permuted Output: [FpBN254(0x0bf747c6db17b67b393a8a8a4a0e3e47dfcdba588001168403e9ba3f827e06fc), FpBN254(0x1f428fac6587d07ee7298d06390e53539b2e6926660605ab4e9544a6d6c4d1f3), FpBN254(0x240b5c1e21e070a3fcdd7cd2a964551d47e54a56847172e639b09e48ff6ceed5)]
 Permuted Output: [FpBN254(0x1f15e76452be89c384650d8e6d0c75b135fe406a1119e99e2086e550bc66b4cd), FpBN254(0x066fe346c642fcc7ab0a66229cce1492e01076753706c2acbb0d9b181494d202), FpBN254(0x26c3d794536367db0d534b0ef74802ba231b693a153c0fede8c9a59690374a9e)]
 Permuted Output: [FpBN254(0x04c971e4fbbf96ca3f12e9af21be4c2d88ee94fe9c15e9ff7a51b7ae4ced5723), FpBN254(0x1570114956e966250b6352009b376ebf524ccc6f865543533148486044c9afef), FpBN254(0x158a5b4f2c41e9fb9ae86307c6c58a20ee19850751d5d1ded0b1148238af9984)]
 Permuted Output: [FpBN254(0x21ec76292069dc6b196a97814fc77e4fa09869399cff347bd0396281ea1d3141), FpBN254(0x1e4620d096c8c28e45afefd87609dc6c5339e9ae3342f60a32030c642ba8c5e0), FpBN254(0x212fb94e1a265aa9b75bb9e4101f12ba11b49ab51af2935602bc2bdfd6d61915)]
 Permuted Output: [FpBN254(0x23a9bba6c60e6ac1489892c51048a67884fbf6ee7cae889d91db83e748935481), FpBN254(0x09991d896814dd54c3211634fe9b03b2e12f3907bb1f5b2856f1fa5ea218fa2e), FpBN254(0x16afbfc998efba58af670eb9aa636d08e18eb74cbe52a5a46379dda68ee835d3)]


 
Input: [FpBN254(0x2a695c68be51e24419d80c945a5f683a9e848a996a494b4b0aab2d7b8f6f5021), FpBN254(0x092a4b0caf633f5b8249a766885a7ba5edb79fa0f229a0fda99047a4ce1c863f), FpBN254(0x17ef829dafac978b16ea501e4cf8d1dcaafda86a6db4065d029a2d248c415cc8)]
 Input: [FpBN254(0x1cdf2364327771226cb1f9f28953747f3c24caeae8dea3a5b9fe22813dfee730), FpBN254(0x29ec3a55e910691fa11422e5d7c204b7ce1d580331df6955e96b85caec76c4b1), FpBN254(0x2ff471376d9b5e5ae880996fb5e3e24795506d6cd58cb7d583cf0534750f11d0)]
 Input: [FpBN254(0x0cc96fa8cf18423e2588ae2ec146fd40185800db2f330486a97818ded2bea32a), FpBN254(0x033f7e91a97fe3f008d05ed0935b3dee5940dcb4eda61b91cb0d1dc7659bcba8), FpBN254(0x1baece0f8567b5a469b919e40e6fad296972289ed698e932b35f694fc1a109a0)]
 Input: [FpBN254(0x2b0d64aed0d40016dcabdc773a633d19f84da10cf39a02a97269a0e85778ba08), FpBN254(0x18b4d6511a2b7abd1c7be551cecf81f386c07945597cad022e0aa3defc88ee9c), FpBN254(0x132101460bb2325a03922e1b5c7d800b34d5003ec3e455b17a9c9ef13dcf6b90)]
 Input: [FpBN254(0x0ca7a1ccb3601d4390d665c78ce05f9456899ee269f09b2fc510a52306dbaa0c), FpBN254(0x1fedbf654acfb7ac5f8bfbe16bd96c97ed5888a07c2b212e5eaaa653ec96f125), FpBN254(0x0c024aac1016eec32f24570df1d5cdf05faa6411333e57a8993451fa78888a00)]
 Input: [FpBN254(0x2b2823586c620a87228a8b28e4a5aac5baf05c4d950636031e98ac7dd874fd7f), FpBN254(0x1d7df4890d1ee9282c05248e92a1dc50e94ab4cd28eb7347e958dc0e6e019782), FpBN254(0x2d2ee35f01d2e7328447df2258f796029bf7f908552f1faab3f4987ed2f166c9)]
 Input: [FpBN254(0x297c8fb92eac1654c6136dc57a8f0be8c54376d87c155c9f06e6e7f5863758e5), FpBN254(0x0f3209371bd8553a6ce025f27ed9dcd14c76eb27671c9f72e88a932c6664cb77), FpBN254(0x16caa9facde5346d6a81c786855d1fa1de0c26e462e6c6a498f61c77c40b2822)]
 Input: [FpBN254(0x02c3013a366483e65169db4c20fbeb86cfceedd3ea870b0f8f69eedf771e6d80), FpBN254(0x070b9257df50ef3af275ae13b23e84ab8d70703e48d13082c977ce07c98c485d), FpBN254(0x1b0350431ea8c032eabbd00429ef0aed7066bf831da98c97eea86c804a1b9f09)]
 Input: [FpBN254(0x0515ebb904e11a223a1a7a117778cfe10e1f8c18dec6eaf7b0f9bbc0855e3311), FpBN254(0x0cd821a004940d9ffe2395d85aef848f9413616027348bc4ef75990169b39c42), FpBN254(0x29849bc40471f4995859aad75767b0ab75a4923f62b719e2f32bb520d25df6c4)]
 Input: [FpBN254(0x0d2c10c0aeb22479f4375ae0c1d72bd094f969c91bc893febf4711c99d9f4d52), FpBN254(0x03226d3e6077f9994b47dbaa520a56d16507564d112c82bb61fdd9d424b712f5), FpBN254(0x2cf8de71836cba4a7cbdbe7b591b00517253becfdcb2fe9fa276650b1fe50ff7)]
 Input: [FpBN254(0x1f9e13f78cce312f2437f9537543f6ea93156e361b5b545b748047e8ced18642), FpBN254(0x0fa287b5ea4cfa49e6dcf4df983436cc72622d45f63f043774015f3b4540d7bc), FpBN254(0x014e4e0d613fed9ba6571ff42d49381c07e58cc38c6f3e90d14af0c55b9598a4)]
 Input: [FpBN254(0x191607022b1d68284cff3a99c1bd77ee757e9a69963924caf0b5599b90e3271f), FpBN254(0x2c5a7a472b5493b29caf8c3a712310b8c24f33dfa87620be56db9b3da42c83d8), FpBN254(0x1ea0d20736a52898695c40fa37341694feb16184fa9aa9293bcd8966f14958dc)]
 Input: [FpBN254(0x1498e7fdd7e5391b73021c322b69aaeca6d5f7f4d8d18c63152f0a928aaebbf7), FpBN254(0x02b717354a832a9e7e070b0a0833f063e006e5ee258bba1b9175d5de73968ccd), FpBN254(0x0cb97579e3d27994886d949abc103062ed4711b44ae6128d7682bb60e9d67ab4)]
 Permuted Output: [FpBN254(0x2f6c05e6495794510f72edc18604a3efb04189d9b5cc2898b92e52748b4226fe), FpBN254(0x20197312ee86c1290a56394d855ed52e62aedf7ac544270b7a18ff05ef780ee3), FpBN254(0x2b04e9849c0e30ef1d959a985befaae21ddadd18ed54fe39f99c8c28e4a1654d)]
 Permuted Output: [FpBN254(0x1e11faf59ce2978c3e7c514a71f537dfac40156dfeba6e7bdc5ea68ac8268e72), FpBN254(0x0ed6327707e7bcfc0188550838c281e49ac52a1b7b23c6369b157cbbe4374539), FpBN254(0x29af37b73d237baf25d8774ecce47224348f68d4ce1e40f87476bb621f839b2e)]
 Permuted Output: [FpBN254(0x1b9bdaf767a0e9ad6302643fec5e5b06605d4d2f062c3c97f153e278b793a851), FpBN254(0x239371153c3a4ab0a928bc82dd88958037e473cccdab58571e9a599dd7e5b9e8), FpBN254(0x03c059312478c67657e61443c14966d98c4c4d6e715ef9699cf5bda9f782396f)]
 Permuted Output: [FpBN254(0x24b92a162757d3c34f46ba816e431935a7e9b5da5f8f3ddbbcf7442bc60acd14), FpBN254(0x1b1912b82d9ed9901df81632fc3e8e5ab770a03dbc8a50aa883f78d3a6dadeb1), FpBN254(0x20cb26a99a99d3302fce5295f9bcf7a525df0250eab640c99901d03eaa5a1eb1)]
 Permuted Output: [FpBN254(0x0fc787d2ebcfb2aa79e0a18166d69b876b9576eeefe73c6e2c5dde1f8466dd7d), FpBN254(0x0cd14557b89e84641a6d6c2abc26df43b992e1e77bfa30ed299035b1329ac80e), FpBN254(0x01c49d22eafe9709ba2576e35301aeb5e1a1efdfa1041c76107219be847af5d7)]
 Permuted Output: [FpBN254(0x30451b7d63f6a8b5790d7e99bba037076fed5fb10c17b97e66d142a2f6e73614), FpBN254(0x28c228126b266c55271b8e4c4b9d9d43cde750a9587e8eb861daa582999d22f3), FpBN254(0x14d98be7535dd85f5c248aa9e223212055aded6cb53f877fd6f4a975ae95bfb6)]
 Permuted Output: [FpBN254(0x20e4272d0b235cf151d0c1afb8d0941380c881927d81a29ea651faabcf437002), FpBN254(0x17d357bf21af0e6e169845707f62fe1ca42ce18655bcaef15f4ef7d2d1991653), FpBN254(0x05798f489212e114bfdcd5b53144b97131af9ca8abd240311654b03068bedb7a)]
 Permuted Output: [FpBN254(0x20b924516a2494a8b6fbf8ade3e7d646c2027eb268edddfcb8cf4a1a137c7b92), FpBN254(0x1a921ca46e7a09ae29d0cb1ee1ac4748716071f656e21bd7c70d47e470373b9b), FpBN254(0x1ad65327b934656c2d7eb4c81bcadcee6c2bbd2796b42844c330a5aab12b8b56)]
 Permuted Output: [FpBN254(0x2a806e61e406ab08bb3b0657576ff81e447f2709553050cff623dd74dad58a49), FpBN254(0x24de4ddf0a229fcb4483cb8d2c8b13bf8f55ea5ab7c3bee09137ea3aa0df1d41), FpBN254(0x0ac9b4cfd451cf9a550cf65ad7501480d7fd3a9163034bb1ab6d5800c59b353c)]
 Permuted Output: [FpBN254(0x045479759d8c625b15a0a553cce88104910328177e71a9cae5ea8c33a219cb93), FpBN254(0x0f27addbd42b1aae3282d5e15c839ef23b71ae1a63296526b298cc30f87571de), FpBN254(0x20d4906bb8463af5bbf9a7ed4f8fa1a4b8bee8126380b736b39aa6fd2736777d)]
 Permuted Output: [FpBN254(0x048349dfed70d26a4e0daa522ca268f865686cb77c8b6a602d32f42a7fe23a90), FpBN254(0x020adec759446020552a7ee308f748cc6cb71638835f583670f1e379ea779beb), FpBN254(0x046f76b6e734fc6017649e41ed6437e4b1490c96e7236d03a4abb5a46798e0f3)]
 Permuted Output: [FpBN254(0x1e1b417647aaadc77c3409dcb552f16612e715ffcdd4fdc23a53129c148a2cdb), FpBN254(0x08feddb39ca46924f43172ccdc7b8ea717277505dfdb094de1984cae14aeb3e6), FpBN254(0x1f293342f446633fc639a0089568c7c116cdeedc3f55891e198558b537f89052)]
 Permuted Output: [FpBN254(0x00746822205e9917521f6f6319965589dfed9caabcf6bbf8917c86c9b8e9333f), FpBN254(0x1744a8d8667c0aaab9d6fb51762aaf71853db37e5e35c61f4605e4ddf8ba4c63), FpBN254(0x084702e55dc7ef84286a1adbcf7bea7e9ea1af977a837b328bbab5d2146a5d32)]


 
Input: [FpBN254(0x014eea4477165c9e5c417d5dc235ac59eb463a6deb1174a608c3aae2712f3586), FpBN254(0x13b6e317c2bd226baffd9ab9ecd6f22121aef3569120a57bce01f2067b96376c), FpBN254(0x0a95bb4044e2405ada9082d84e894d2ed9f3e1a6ec209a54a2a91e416ef7dc55)]
 Input: [FpBN254(0x10961d47b26d487a4ff9b92aab1bdf78d7119b3e88196d10f9d9e7fe6098a285), FpBN254(0x1e2dfeb3f6615d2b91d8e4eaccc67bdc556eedce87494bf92020121ef8f9ef57), FpBN254(0x045ec3f0cff07b3efcebcf8fb0808c31349affc96a7c07e32865f8a08d878020)]
 Input: [FpBN254(0x01d97a55d7354602f331725ad35f23f269c184ade60a03e349e0d22e9eb1ed00), FpBN254(0x01914c5505542f9239bdf67c2d7fe4a83adffd8e01eb54b50bb227ec248fd9a4), FpBN254(0x24e2f6600b83f0e2ac818524639e34e4dadebee6f3dcb6a5f8c2dd579c070b3c)]
 Input: [FpBN254(0x2f42128a34b5e0848927aad4c1ddf2cacd0e433bb6049818c633bcfc871d22b0), FpBN254(0x0f7a1132c92c780218970d3e8db75d05c6b7e6d7f45ee5c09b53fd445a788414), FpBN254(0x1ce1cae19ebb796f6339ea9efc152e5a827ac0d032a7c9d4f8582227818dfa9c)]
 Input: [FpBN254(0x2dac405dec1c57c8ae85b5bd4cbc75179ffd20a78a8ec6770949f1a030b2f7ba), FpBN254(0x2b90bcbe97afa8391fdce131d73ed74a6bb6b5a2c7b4a50df7d91ba8493eed67), FpBN254(0x2f4d851ab1237715e66cb242badd36765681d5a3c9898b4f4b33d6863f287c70)]
 Input: [FpBN254(0x305ab23c7341d81a5b905e8966c80c1a6e7798060e506d88da161c2b4c957906), FpBN254(0x2730939da1381beddb260cd1aabd7c9b0a766f383fa68f7ccb688e275f5e4ed4), FpBN254(0x108c6af7950c938b182cc3907e361bf6d88c7407c797595821f2ddfced6a55c2)]
 Input: [FpBN254(0x0dd37612425c662c8251ff379eb5f81ade4dda5c6b113d5bc86d9c99d285b63a), FpBN254(0x129df9931c75ed619af24982397c03aff096202d1b840dcf865ea93bd4c8b15e), FpBN254(0x29dc9a6c253d6c43775aebc421414a3938270ef012f6a05e4695e4622055bd9c)]
 Input: [FpBN254(0x006690d52ff3c403a8b5f948946dba308874e955e6d6d6a77f894645487e8668), FpBN254(0x058212eb91f6ac1e5856a457376c51e9adeb5901f1dc007d92f3b5e66bda030f), FpBN254(0x0e45eac734a0f8690c603f1f2bcb0ee3c8a050247248fecea68267dabc7a7bb3)]
 Input: [FpBN254(0x05057bc4bea006bba8784caf82a5f9276caa050ec008d715ca1fa0f0c414a1f8), FpBN254(0x1800f4844426741e726f2f35e38b6dce845946711326a3c3abd4f425629e4702), FpBN254(0x12c8aef69538ef45be8beb281cd6057196ef1468f9317e92ef6298b6f7cc1993)]
 Input: [FpBN254(0x02f1daff38e4bd57401ed88cfcf857406a16d82947a7bd855dfad33bbb74a6f5), FpBN254(0x18baa64f6ba04fa6c1864e03e3a3e591afb4550d795b0cab154b17d05deda1aa), FpBN254(0x1d1b4989d413488ac4c3b17120aab25a88c250b03a2441264de194ece64b8ff9)]
 Input: [FpBN254(0x1e86f19a7f26a73b99f41773cbff7ca050a59e8e135af2323bacd5e3c19a0a98), FpBN254(0x08fb3b8504f6f23f66dac82a6ed9af7927b8cb1ef8d927315c5f03ef76fd82f4), FpBN254(0x2140a8b2913fafaad3dcf80e499f4965c7555d436f92f30fe78edfd424183797)]
 Input: [FpBN254(0x2060925074428762d74d15ea32fadb16717e4ec359c340a4ced740f300c48c15), FpBN254(0x042429c26d815dd3aad1763cc7edb5f062b9a681b37196734a9edf3ca6758741), FpBN254(0x2f72ce231766dc44399f09a6874b73bbff782d48c1730c073ac72ce0046a86ad)]
 Input: [FpBN254(0x125003f72b6f76a8bc227ad80de95f19de807904ff1155a892aef83b17ca5f2c), FpBN254(0x12e073dcd8154d8edd5c5b3d5de8c42deb810365d0b2a0bce8a4d263d7f973f1), FpBN254(0x180361c198fa2924e65c831463c1ef80b8d07398d433c37fbf77ac378426a25b)]
 Permuted Output: [FpBN254(0x275b5d6131dad6693281cc5c982cd5c8511fbcdb10dfc7773d2d8507a7ed127b), FpBN254(0x27082dfd11395f0d816f1bbd2c8cb02e075c0a2b13192b88b0a0eab05adbc193), FpBN254(0x1314b4a1a2162923c293a7ba482c066804c8771da591aa533f78de24759905d7)]
 Permuted Output: [FpBN254(0x1a3028c87f475c359e0146d51ef97acd875329cff23f042e86e010a5c90bba25), FpBN254(0x00756fd99f30cfc7cca85ac478074d63b8f0b92d355e94bbb533d010f2f9c042), FpBN254(0x2992a4e70f533a804a327dd2c85798ce3576eff7b9019b810f7f193b23e1e88e)]
 Permuted Output: [FpBN254(0x07cc376892cc5bd0a0b21eaa4688e1e69ce3b8f13873384911e155acaeec934d), FpBN254(0x2856befbbf0752a37e56583cbb5639a2be33b93a4eb0dc81b8a1876526816930), FpBN254(0x164d360a6f4bf510d1c0ed77c6aa9a41edb8fd25001f9cb4940767039ca2749e)]
 Permuted Output: [FpBN254(0x08b1d236eee421da956e384d228a229c6b03bffb8577db443f8e5c482ec3c088), FpBN254(0x29fad7d77c54acf872ddf1d704d2bd5ef220675761c3787621c1233e9c8d3e18), FpBN254(0x2151a4d4f2ff7335620104836a413c549fb029513a94addeb55a860dbb7b98a2)]
 Permuted Output: [FpBN254(0x0b443c1c1414b1f9e2e4f14b28cbc1569701dd6911dac1ba080f621b8529ddb7), FpBN254(0x2aaa3e566e2725392b46b0f359afb305965867757ec5adf2354ffc056567f0f8), FpBN254(0x05b7ed78d0cdf13f9a9ba87de6c9d88e45617acbf6431c0fe981721e8d9d7861)]
 Permuted Output: [FpBN254(0x1caecf120390a1e4d6f6ef02095d722025c4a24bf781d4a700c21bebc78a9d7a), FpBN254(0x21deee39f2eff549ea0d85b749b7db58c95089e1bb196eda0b0e8e7a73e77064), FpBN254(0x24ac53dc2b42ebefc59c939d023354bb506c501ea786fa0197117bdd78d2e15f)]
 Permuted Output: [FpBN254(0x023dccf6f7c6e1f7902b68c0f5217d6d8f01f4982237a307c674e1ce64e9e4c5), FpBN254(0x246d1877b9d608943202aa86401e163e21dd41b41cda4c88ffca36e71dcc1ed5), FpBN254(0x28d272cbeeec71cfe0d961980959fbe7c5e6af089c29a110301bfeb299b4b201)]
 Permuted Output: [FpBN254(0x162c413c452efb0bf617e3082b53b03864464a430f2e3ed0719a15c21a968339), FpBN254(0x04e359461a33bd45d55cdbac35d42a829920e7d8016d84df684d070d5a547eaf), FpBN254(0x0f00a8c035a24e3367e8596b56cbd84efef3b3742522c3d45549f9b292112f32)]
 Permuted Output: [FpBN254(0x2ac31b4618ee4869be90f827860b7d90bc8f5013271487efed3b43656e3e47ae), FpBN254(0x29e31f576bd333ba533637b022cbcdaa2380ffe5a75f1bbc915bfa90c2c210d0), FpBN254(0x27be15feb0a84e24f2f8edde7a7e8b99542407fb728d7df0855506d47c314424)]
 Permuted Output: [FpBN254(0x26e8e8839b22cf312112cf59cd789c52a277d1805fdf14f66152b6dfc68ccf8f), FpBN254(0x0d1d80746e2bb726b3ae572e34fd0bb371970fc741c590b618bc219ab3a59ba9), FpBN254(0x27c11370de75b4c9ed85f348e716d1d7ec89cdf3601353e93cb17370fe3a2417)]
 Permuted Output: [FpBN254(0x0638e5f31432db876cc22fe520d2e20c10b0c6b26c296d467e9a0c431604b616), FpBN254(0x1b1aa2222e531219f65f2f1329eaa67589fe22cf8e348999a4d2c268c7e476b4), FpBN254(0x1ddd83d8282cad70f571a7549072c84609a0f573e9af080f08015e05b9131b20)]
 Permuted Output: [FpBN254(0x16636938b4a4367ccfba2f75e282c7ae09c250884a3136b5da6fe9686460d27c), FpBN254(0x0ff87f08e3e124692875b3c3c769ba35e11ad64ee8b3bc561de5d23a1d7e2411), FpBN254(0x054f358a986362487776e6f3fef08b3fa05fe95b62e319fd046f47b9f62f3190)]
 Permuted Output: [FpBN254(0x2113e97a98ecf7fc1d78406b98e819557b18da172d10d5663b7b72895af693bf), FpBN254(0x18dce19f415518ce2aeba590543c9ded9cfee64e27d71117c499af8310617de5), FpBN254(0x17bb6a91791a56b169df7f9bee90b990946cbe863417a081fd22e4c2a22bf576)]
*/
module testbench_griffin_v2;

    // Parameters
    parameter N_BITS = 254;
    parameter PRIME_MODULUS = 254'h30644e72e131a029b85045b68181585d2833e84879b9709143e1f593f0000001;
    parameter BARRETT_R = 255'h54a47462623a04a7ab074a58680730147144852009e880ae620703a6be1de925;
    parameter STATE_SIZE = 3;
    parameter NUM_ROUNDS = 14;

    // Inputs
    reg clk;
    reg reset;
    reg enable;
    reg [N_BITS-1:0] inState1[STATE_SIZE][13];
    reg [N_BITS-1:0] inState2[STATE_SIZE][13];
    reg [N_BITS-1:0] inState3[STATE_SIZE][13];

    // Outputs
    wire [N_BITS-1:0] outState1[STATE_SIZE][13];
    wire [N_BITS-1:0] outState2[STATE_SIZE][13];
    wire [N_BITS-1:0] outState3[STATE_SIZE][13];
    wire done;
  reg [N_BITS-1:0] testVector_1[STATE_SIZE*13];
  reg [N_BITS-1:0] testVector_2[STATE_SIZE*13];
  reg [N_BITS-1:0] testVector_3[STATE_SIZE*13];
    // Instntiate the module under test
    griffin_v2 #(
        .N_BITS(N_BITS),
        .PRIME_MODULUS(PRIME_MODULUS),
        .BARRETT_R(BARRETT_R),
        .STATE_SIZE(STATE_SIZE),
        .NUM_ROUNDS(NUM_ROUNDS)
    ) dut (
        .clk(clk),
        .reset(reset),
        .enable(enable),
        .inState1(inState1),
        .inState2(inState2),
        .inState3(inState3),
        .outState1(outState1),
        .outState2(outState2),
        .outState3(outState3),
        .done(done)
    );

    // Clock generation
    initial begin
        clk = 0;
        forever #5 clk = ~clk; // 10 ns clock period
    end

    // Initialize inputs and run the test
    initial begin
        // Initialize inputs
        reset = 1;
        enable = 0;
testVector_1[0] = 254'd21522355681653392990718421087354924920017962571854039821646797661308615193169;
testVector_1[1] = 254'd12474386525783842807182291508500613291262455221924536584473603971436929495095;
testVector_1[2] = 254'd10854212365580904016637868862894703901217599761197551470531703969797269735423;
testVector_1[3] = 254'd2833974035242175361896882010450368535794379467427702350262701998395342954978;
testVector_1[4] = 254'd13768265560189264423348624617942974097115584620159875324125610057825582650234;
testVector_1[5] = 254'd19475427961875606093009944485797249498742278763348943538250751354183624528287;
testVector_1[6] = 254'd16077998017997257624383264093330711462905255408438113761799522589399789066424;
testVector_1[7] = 254'd4591336034794362249429651446012613609421789048335211440180260414985675979571;
testVector_1[8] = 254'd9581701609975595081371886836405626672681585559807644047120794916609717516335;
testVector_1[9] = 254'd9934228559362985316616133250034310015267948255228817288726841870317183643433;
testVector_1[10] = 254'd3913437246589357335193816422522758473852965250950193924635313438966189344627;
testVector_1[11] = 254'd5845552450062575214067131224394954485922860972448369992559201456849681162227;
testVector_1[12] = 254'd4774618147654992938654428650511445935175121931017412153575385320392655695810;
testVector_1[13] = 254'd6608546553117878864031299337550523869901158948493997119628170326836658585899;
testVector_1[14] = 254'd2476114185100296265626846695706034421507349737697405629650360613089094646953;
testVector_1[15] = 254'd5808003784028367785172025847890330892647915296548678014622262346567814302080;
testVector_1[16] = 254'd19409774051401924034233771314033459553278905591721948434108726533191567834935;
testVector_1[17] = 254'd7275749124359065717739904581567875812241985553742970107527303279095757564628;
testVector_1[18] = 254'd6833700902594805773105324002200552098484020285658907442900270070294614862521;
testVector_1[19] = 254'd17508011390153325253271810550118415735250948930242972186128259135103397854820;
testVector_1[20] = 254'd6186010267483752614335520235028749204874024605643955590546498061892261214341;
testVector_1[21] = 254'd6256977619560381777693174096563571844113964742681044195644485266580221141912;
testVector_1[22] = 254'd2564144855453765267488568411854410167500670465814170043330172684818008191346;
testVector_1[23] = 254'd8901823469592236431327715215262749442802410294294994492863032136604209717096;
testVector_1[24] = 254'd18813502421346713446774187286043312846165805210826842266475429766958069832730;
testVector_1[25] = 254'd3382234311100456351427862291847096994612876427512386703811661003015106691317;
testVector_1[26] = 254'd5172685326803830614001662263565268020658487588553384094623727583751542007216;
testVector_1[27] = 254'd4295172293365356772888468616978025967128812415910130942968508160521997459667;
testVector_1[28] = 254'd10481398846165754052582941953393973996877778032366087850394796618312571882170;
testVector_1[29] = 254'd1771818477988466772902754635620828869424254897413195973088354838058158723872;
testVector_1[30] = 254'd2956326865233873909159814639276832934954702793571210378275049393719348936921;
testVector_1[31] = 254'd18477027113244290334479136841868667171247363331452115693114275427050144601129;
testVector_1[32] = 254'd17612464637965053291913205295942475169085498897537073614858704702365730275835;
testVector_1[33] = 254'd13466824521569867727471394352850610930668768478397876229032222252136220495003;
testVector_1[34] = 254'd11006050214562741459871684086456412916114677564947055823541467039134264012534;
testVector_1[35] = 254'd6077301026332713992608446293548860164795750449247318481245176826584014837193;
testVector_1[36] = 254'd12256044551403186078225307486729203329869149386393174200336715764728961844772;
testVector_1[37] = 254'd9293384229337912360401493586773195282365182255236744587766889132141157990592;
testVector_1[38] = 254'd13346508422652734171563656901046034884051028058908505815988821769554849589383;
testVector_2[0] = 254'd19183296366840297261607075654228646741064326077950506146152119958439979864097;
testVector_2[1] = 254'd4145541186935938026593050205566893848843983243153598113321915732773859788351;
testVector_2[2] = 254'd10826373444134521561985703079771848275272288331843813040865871873516991765704;
testVector_2[3] = 254'd13059010918208593108840516037810737021500968883900878897087531485752054441776;
testVector_2[4] = 254'd18962205316629716089629550045781349996410263508838025262691497606025043166385;
testVector_2[5] = 254'd21690595958896654773242916386694403137299006628807566917516254018927139426768;
testVector_2[6] = 254'd5783661087944809595360845793696567520915671280836123294983292365757143229226;
testVector_2[7] = 254'd1469123457913188069101400702126786136560629096678798972410169925466448448424;
testVector_2[8] = 254'd12521300479215468644919198612302506167495523179877046350617389170802716379552;
testVector_2[9] = 254'd19473116388580141389032591771207874584755915878881382939147643628206069168648;
testVector_2[10] = 254'd11175019997888401711022850064888905062154712112269322475742785655155102117532;
testVector_2[11] = 254'd8652258866394102626161833837856845832809035066075201407074359983062031231888;
testVector_2[12] = 254'd5723934342698579566388545792479377786322174066748665471581872922956987607564;
testVector_2[13] = 254'd14441762024819145101563312900197271935433757243634442358857277566865458524453;
testVector_2[14] = 254'd5431803245163673298976842365073723058211043027681474475943116161740421237248;
testVector_2[15] = 254'd19520370316683093731719802927983557890256086175586465383333423001067383487871;
testVector_2[16] = 254'd13339616213015109345825002458705833605132322667027309331536391930989519148930;
testVector_2[17] = 254'd20436922409034520793965692692214297806629627496041500534582526246916461782729;
testVector_2[18] = 254'd18764907770179324051153353341835142085078612376154171345987645895951097747685;
testVector_2[19] = 254'd6873098683434528928059976161039078516855136952707773929571866369873510976375;
testVector_2[20] = 254'd10308958932719677747283778537406565112470406926683357228987760894100332292130;
testVector_2[21] = 254'd1249169345949784524964855429711449940529535943731343235391962195486771670400;
testVector_2[22] = 254'd3186635281795353972101562547598207898460383479097088651952210749978632276061;
testVector_2[23] = 254'd12218301402195486376443806165731614872580552908260829499993774131958041517833;
testVector_2[24] = 254'd2300294929772158011405127391373343360703354444240793700720222120249982333713;
testVector_2[25] = 254'd5809625220694393238157569615612389671746093850556705662627995764004041759810;
testVector_2[26] = 254'd18779125659766095679587997652319628327081884848497819919219193669738859198148;
testVector_2[27] = 254'd5957923925081643019715130710860620413793722037983904528875544661238317272402;
testVector_2[28] = 254'd1417765317980092617695561343387852538338397354720835260057582354060035953397;
testVector_2[29] = 254'd20341478657732359485015097777465126710742012188813049535518454386625878495223;
testVector_2[30] = 254'd14300997949432201924743277685599246443944405833844689704363257305644364039746;
testVector_2[31] = 254'd7071858593425000602801186179750089534735017278159141702530112743926480820156;
testVector_2[32] = 254'd590665616571927512988326133754589685197369799085150979574811949155772373156;
testVector_2[33] = 254'd11346740220691630857148898955135667519757521554470402151610280345499670357791;
testVector_2[34] = 254'd20061625505267518973076494615914930073089394071518635780390141135042462385112;
testVector_2[35] = 254'd13853530549069791879699142905485692307325268623244667738444995055667273881820;
testVector_2[36] = 254'd9316418872520697207326607613630008938336898439318906321463318135026215730167;
testVector_2[37] = 254'd1228118886911194995007031869401821156972588644036210345341629112411777043661;
testVector_2[38] = 254'd5755431680451793552524807876072280996525815020491463183965467442175681133236;
testVector_3[0] = 254'd591743774098864540218411108332085793609522769830409381750210192903662155142;
testVector_3[1] = 254'd8917077625879612115413971842737879523287250565580797868493049778358174758764;
testVector_3[2] = 254'd4787681057742389937194061545882083283900123257827609584518295732975962676309;
testVector_3[3] = 254'd7502234720639834540952715783372213958364418729978988072927067674806278726277;
testVector_3[4] = 254'd13650651470762434123907266741255318507155839663563956184860025153971736407895;
testVector_3[5] = 254'd1976687351245630654158196769008656986547990305338716805606060735005389717536;
testVector_3[6] = 254'd836562988954009092784030740652587056070884621420094368982282415366261042432;
testVector_3[7] = 254'd709032497855148404822425443172153488055950547218216665850808674287625427364;
testVector_3[8] = 254'd16684270404606407935670470434755543737013503676595466570535495208689037937468;
testVector_3[9] = 254'd21375443747146834950281329619159540790843387873838572513280231381248006496944;
testVector_3[10] = 254'd7000366769523251532158389334154541546608156937511165619596891087487358239764;
testVector_3[11] = 254'd13063700585373111711769804124488051749810544890634396199199266858628423744156;
testVector_3[12] = 254'd20658420125295464651570027671343501486913149935527574106807264182660991481786;
testVector_3[13] = 254'd19705181133086022618628978689550110324431098896255788148274315820660867132775;
testVector_3[14] = 254'd21395669759279057491132093412251347028818447829707472228479349082473336700016;
testVector_3[15] = 254'd21871263108411370235982499998915474761683948113640352479861461458528199080198;
testVector_3[16] = 254'd17726028560259717452720860269887091878272601877840500674346010755921176579796;
testVector_3[17] = 254'd7485102426317527671373743126224905929296165474723370424706359392066463225282;
testVector_3[18] = 254'd6253686660587285479645320767173657882033235822713528960121162830555921102394;
testVector_3[19] = 254'd8420748764618768884007413389394142756417758336635926082733054446391593054558;
testVector_3[20] = 254'd18934598930698634983943919344033433353654851627182383078629747610201651264924;
testVector_3[21] = 254'd181217999599930238993371861800689473097957051209352083640365424785848436328;
testVector_3[22] = 254'd2491384943730988321299738271343162216888943199113909940621891291025220698895;
testVector_3[23] = 254'd6455912706852432239963302770735825870908835943080032306559086820804274060211;
testVector_3[24] = 254'd2271252697265592283281665725590763527281049768366349219051950182687820784120;
testVector_3[25] = 254'd10857195957997025005096914296272638114081102168013591485009484765336273045250;
testVector_3[26] = 254'd8496208239180646552195200843921249194880206562995078385304811537846332299667;
testVector_3[27] = 254'd1331947301259710218671988446450552570460347260048775200383407567904219375349;
testVector_3[28] = 254'd11185289751110890130429592949951618081159123751242889404082324494237844742570;
testVector_3[29] = 254'd13165285022993889301504559418373242013825165698144166210851981969271089238009;
testVector_3[30] = 254'd13807810450270220486413823048511392044614673759083339713584365222972150647448;
testVector_3[31] = 254'd4062392191155709921946143084245794572981995459228520722542094612326124454644;
testVector_3[32] = 254'd15040566522946856256121711789780703993906044174915705088993624123250887374743;
testVector_3[33] = 254'd14644638296889208333770065316794673289389943045135246880216745076247123758101;
testVector_3[34] = 254'd1873146102027217317439075170827330600958025652568975468817846258402359347009;
testVector_3[35] = 254'd21461547154608325302745365567747108938063852689921886788689379285405608347309;
testVector_3[36] = 254'd8283006408601214866054875973330118908400529610020209611015986704865261412140;
testVector_3[37] = 254'd8538204671783519298862696591580388040565229941315494469410659783235969053681;
testVector_3[38] = 254'd10861483595968452403246580609824210412656714897278200188349520796347739316827;

        // Apply reset
        #10 reset = 0;
        enable = 1;
      for (int i = 0; i < 13; i++) begin
        for(int j = 0; j < STATE_SIZE;j++) begin
          inState1[j][i] = testVector_1[i*3+j];
          inState2[j][i] = testVector_2[i*3+j];
          inState3[j][i] = testVector_3[i*3+j];
        end
      end
        // Wait for computation to complete
        wait (done);

        // Finish simulation
        $finish;
    end

endmodule

